library IEEE;
use IEEE.std_logic_1164.all;



entity DecisionTree_tb is
end DecisionTree_tb;



architecture test of DecisionTree_tb is
begin
end test;