library IEEE;
use IEEE.std_logic_1164.all;



entity Node_tb is
end Node_tb;



architecture test of Node_tb is
begin
end test;