library IEEE;
use IEEE.std_logic_1164.all;



package rf_types is

	type std_logic_matrix is array (natural range <>) of std_logic_vector;

end rf_types;
