library IEEE;
use IEEE.std_logic_1164.all;



entity DecisionTreeMemory_tb is
end DecisionTreeMemory_tb;



architecture test of DecisionTreeMemory_tb is
begin
end test;