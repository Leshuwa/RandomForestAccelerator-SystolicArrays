library IEEE;
use IEEE.std_logic_1164.all;



entity MajorityVote_tb is
end MajorityVote_tb;



architecture test of MajorityVote_tb is
begin
end test;