library IEEE;
use IEEE.std_logic_1164.all;



entity Comparator_tb is
end Comparator_tb;



architecture test of Comparator_tb is
begin
end test;